library verilog;
use verilog.vl_types.all;
entity Disp_VGA_vlg_vec_tst is
end Disp_VGA_vlg_vec_tst;
